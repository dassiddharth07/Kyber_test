`timescale 1ns / 1ps

`define     WIDTH   13          // Word size of coefficients
`define     PRIME   7681
`define     CONST   8736